
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h4d12822a;
    ram_cell[       1] = 32'h0;  // 32'h7efc6cc6;
    ram_cell[       2] = 32'h0;  // 32'h7023e40c;
    ram_cell[       3] = 32'h0;  // 32'h37eb376d;
    ram_cell[       4] = 32'h0;  // 32'h9d907463;
    ram_cell[       5] = 32'h0;  // 32'h86ff4f8e;
    ram_cell[       6] = 32'h0;  // 32'h5ac011fa;
    ram_cell[       7] = 32'h0;  // 32'hd2a8b63f;
    ram_cell[       8] = 32'h0;  // 32'h0ab7d6c6;
    ram_cell[       9] = 32'h0;  // 32'h57ce62ca;
    ram_cell[      10] = 32'h0;  // 32'h4cc71bee;
    ram_cell[      11] = 32'h0;  // 32'h844bb59a;
    ram_cell[      12] = 32'h0;  // 32'hf3769cce;
    ram_cell[      13] = 32'h0;  // 32'h0d402873;
    ram_cell[      14] = 32'h0;  // 32'hf660b17f;
    ram_cell[      15] = 32'h0;  // 32'h453f7d7e;
    ram_cell[      16] = 32'h0;  // 32'h7eca0d4c;
    ram_cell[      17] = 32'h0;  // 32'h9ba95bae;
    ram_cell[      18] = 32'h0;  // 32'h9cebcf87;
    ram_cell[      19] = 32'h0;  // 32'h9a18d747;
    ram_cell[      20] = 32'h0;  // 32'hc404d341;
    ram_cell[      21] = 32'h0;  // 32'h255e8bad;
    ram_cell[      22] = 32'h0;  // 32'hf6234242;
    ram_cell[      23] = 32'h0;  // 32'h577ff729;
    ram_cell[      24] = 32'h0;  // 32'h08c0ba15;
    ram_cell[      25] = 32'h0;  // 32'h1479f6b6;
    ram_cell[      26] = 32'h0;  // 32'h926fa367;
    ram_cell[      27] = 32'h0;  // 32'ha06cbe66;
    ram_cell[      28] = 32'h0;  // 32'h158a5a66;
    ram_cell[      29] = 32'h0;  // 32'h010b2d3f;
    ram_cell[      30] = 32'h0;  // 32'h4bc8a530;
    ram_cell[      31] = 32'h0;  // 32'heeb5540e;
    ram_cell[      32] = 32'h0;  // 32'h5b4988f5;
    ram_cell[      33] = 32'h0;  // 32'h7cf8245e;
    ram_cell[      34] = 32'h0;  // 32'hf5ad1ea2;
    ram_cell[      35] = 32'h0;  // 32'h42eb7871;
    ram_cell[      36] = 32'h0;  // 32'h5ace0809;
    ram_cell[      37] = 32'h0;  // 32'h8bc0e15b;
    ram_cell[      38] = 32'h0;  // 32'h46e5f35d;
    ram_cell[      39] = 32'h0;  // 32'h768590bd;
    ram_cell[      40] = 32'h0;  // 32'h40a29c9a;
    ram_cell[      41] = 32'h0;  // 32'h573ae537;
    ram_cell[      42] = 32'h0;  // 32'hded99632;
    ram_cell[      43] = 32'h0;  // 32'h0397bdfd;
    ram_cell[      44] = 32'h0;  // 32'hf636710b;
    ram_cell[      45] = 32'h0;  // 32'h112c471d;
    ram_cell[      46] = 32'h0;  // 32'hbf035146;
    ram_cell[      47] = 32'h0;  // 32'h3ff163db;
    ram_cell[      48] = 32'h0;  // 32'hf90802ec;
    ram_cell[      49] = 32'h0;  // 32'heba4d049;
    ram_cell[      50] = 32'h0;  // 32'h42bcd710;
    ram_cell[      51] = 32'h0;  // 32'h20469a35;
    ram_cell[      52] = 32'h0;  // 32'h87730617;
    ram_cell[      53] = 32'h0;  // 32'h9eb089b4;
    ram_cell[      54] = 32'h0;  // 32'h0679d56b;
    ram_cell[      55] = 32'h0;  // 32'h2428df30;
    ram_cell[      56] = 32'h0;  // 32'h4931a0b0;
    ram_cell[      57] = 32'h0;  // 32'he91f2474;
    ram_cell[      58] = 32'h0;  // 32'h6bb28335;
    ram_cell[      59] = 32'h0;  // 32'h7c1217c2;
    ram_cell[      60] = 32'h0;  // 32'h19ea7d34;
    ram_cell[      61] = 32'h0;  // 32'h0f242450;
    ram_cell[      62] = 32'h0;  // 32'ha1b6ef3c;
    ram_cell[      63] = 32'h0;  // 32'h474520ff;
    ram_cell[      64] = 32'h0;  // 32'ha2ad138e;
    ram_cell[      65] = 32'h0;  // 32'hecb6eb6d;
    ram_cell[      66] = 32'h0;  // 32'ha295ba86;
    ram_cell[      67] = 32'h0;  // 32'h8a613724;
    ram_cell[      68] = 32'h0;  // 32'h6724dc90;
    ram_cell[      69] = 32'h0;  // 32'ha9502afd;
    ram_cell[      70] = 32'h0;  // 32'hbaba5090;
    ram_cell[      71] = 32'h0;  // 32'h2f27023e;
    ram_cell[      72] = 32'h0;  // 32'hf0254bbe;
    ram_cell[      73] = 32'h0;  // 32'hbf86e454;
    ram_cell[      74] = 32'h0;  // 32'h2b2f85df;
    ram_cell[      75] = 32'h0;  // 32'hcac29242;
    ram_cell[      76] = 32'h0;  // 32'h30470036;
    ram_cell[      77] = 32'h0;  // 32'h18136b81;
    ram_cell[      78] = 32'h0;  // 32'h44df9456;
    ram_cell[      79] = 32'h0;  // 32'h9d6c088f;
    ram_cell[      80] = 32'h0;  // 32'h04b3039b;
    ram_cell[      81] = 32'h0;  // 32'h2f7b1e0e;
    ram_cell[      82] = 32'h0;  // 32'h87f04c4e;
    ram_cell[      83] = 32'h0;  // 32'h7af2ad9f;
    ram_cell[      84] = 32'h0;  // 32'hf6d44d82;
    ram_cell[      85] = 32'h0;  // 32'hd4d4cd00;
    ram_cell[      86] = 32'h0;  // 32'h16509818;
    ram_cell[      87] = 32'h0;  // 32'hf6ef2b1e;
    ram_cell[      88] = 32'h0;  // 32'h7976ebda;
    ram_cell[      89] = 32'h0;  // 32'h65543736;
    ram_cell[      90] = 32'h0;  // 32'h2228e37c;
    ram_cell[      91] = 32'h0;  // 32'h25d09f31;
    ram_cell[      92] = 32'h0;  // 32'h4d4c3521;
    ram_cell[      93] = 32'h0;  // 32'h5fc62d40;
    ram_cell[      94] = 32'h0;  // 32'h7fd2632a;
    ram_cell[      95] = 32'h0;  // 32'haea27712;
    ram_cell[      96] = 32'h0;  // 32'heb7b736b;
    ram_cell[      97] = 32'h0;  // 32'h8f60f2c7;
    ram_cell[      98] = 32'h0;  // 32'h51a80db8;
    ram_cell[      99] = 32'h0;  // 32'hcf874b99;
    ram_cell[     100] = 32'h0;  // 32'h3f03740b;
    ram_cell[     101] = 32'h0;  // 32'he765acdc;
    ram_cell[     102] = 32'h0;  // 32'h00b5a84d;
    ram_cell[     103] = 32'h0;  // 32'h35b74289;
    ram_cell[     104] = 32'h0;  // 32'h31db8547;
    ram_cell[     105] = 32'h0;  // 32'h247a3c21;
    ram_cell[     106] = 32'h0;  // 32'h12fc55d0;
    ram_cell[     107] = 32'h0;  // 32'h3c926516;
    ram_cell[     108] = 32'h0;  // 32'h410ac7e7;
    ram_cell[     109] = 32'h0;  // 32'hd1c7ed55;
    ram_cell[     110] = 32'h0;  // 32'h98a126eb;
    ram_cell[     111] = 32'h0;  // 32'hc6c58705;
    ram_cell[     112] = 32'h0;  // 32'h89883357;
    ram_cell[     113] = 32'h0;  // 32'h193f1586;
    ram_cell[     114] = 32'h0;  // 32'h5df6929d;
    ram_cell[     115] = 32'h0;  // 32'hc20969cc;
    ram_cell[     116] = 32'h0;  // 32'hddb1fa18;
    ram_cell[     117] = 32'h0;  // 32'hd3002322;
    ram_cell[     118] = 32'h0;  // 32'h012a24b7;
    ram_cell[     119] = 32'h0;  // 32'h74cdbee9;
    ram_cell[     120] = 32'h0;  // 32'hf5fbc5be;
    ram_cell[     121] = 32'h0;  // 32'h0c289b7b;
    ram_cell[     122] = 32'h0;  // 32'h5c73909c;
    ram_cell[     123] = 32'h0;  // 32'hc820b75f;
    ram_cell[     124] = 32'h0;  // 32'h79c57260;
    ram_cell[     125] = 32'h0;  // 32'h1e3788ba;
    ram_cell[     126] = 32'h0;  // 32'he8caa61e;
    ram_cell[     127] = 32'h0;  // 32'h32616835;
    ram_cell[     128] = 32'h0;  // 32'hfe3f900a;
    ram_cell[     129] = 32'h0;  // 32'hec126346;
    ram_cell[     130] = 32'h0;  // 32'h80bc2011;
    ram_cell[     131] = 32'h0;  // 32'hbab5d481;
    ram_cell[     132] = 32'h0;  // 32'he59adf32;
    ram_cell[     133] = 32'h0;  // 32'hffe6a68e;
    ram_cell[     134] = 32'h0;  // 32'h92914db5;
    ram_cell[     135] = 32'h0;  // 32'hbd32d0b7;
    ram_cell[     136] = 32'h0;  // 32'heafb14b4;
    ram_cell[     137] = 32'h0;  // 32'h2653106e;
    ram_cell[     138] = 32'h0;  // 32'h998e4ff1;
    ram_cell[     139] = 32'h0;  // 32'h7676903a;
    ram_cell[     140] = 32'h0;  // 32'hff6910b8;
    ram_cell[     141] = 32'h0;  // 32'h4b538847;
    ram_cell[     142] = 32'h0;  // 32'hb9f36e80;
    ram_cell[     143] = 32'h0;  // 32'h1bde6308;
    ram_cell[     144] = 32'h0;  // 32'hacfc19f5;
    ram_cell[     145] = 32'h0;  // 32'h563f75f1;
    ram_cell[     146] = 32'h0;  // 32'h0fadbb22;
    ram_cell[     147] = 32'h0;  // 32'h1ab00a3f;
    ram_cell[     148] = 32'h0;  // 32'hefa2a846;
    ram_cell[     149] = 32'h0;  // 32'ha864ba7e;
    ram_cell[     150] = 32'h0;  // 32'h06f5ba29;
    ram_cell[     151] = 32'h0;  // 32'hef0a55d0;
    ram_cell[     152] = 32'h0;  // 32'he63bb47a;
    ram_cell[     153] = 32'h0;  // 32'h57cd258a;
    ram_cell[     154] = 32'h0;  // 32'h71a345a7;
    ram_cell[     155] = 32'h0;  // 32'he41eb033;
    ram_cell[     156] = 32'h0;  // 32'h5349040e;
    ram_cell[     157] = 32'h0;  // 32'h303796f5;
    ram_cell[     158] = 32'h0;  // 32'h27a14851;
    ram_cell[     159] = 32'h0;  // 32'ha4c50b72;
    ram_cell[     160] = 32'h0;  // 32'h02f78f81;
    ram_cell[     161] = 32'h0;  // 32'h98234556;
    ram_cell[     162] = 32'h0;  // 32'h57a08fbe;
    ram_cell[     163] = 32'h0;  // 32'h05925e8e;
    ram_cell[     164] = 32'h0;  // 32'hb031d0de;
    ram_cell[     165] = 32'h0;  // 32'h6efc5ba0;
    ram_cell[     166] = 32'h0;  // 32'hb48d319e;
    ram_cell[     167] = 32'h0;  // 32'h3ab00a39;
    ram_cell[     168] = 32'h0;  // 32'h2ad38b2c;
    ram_cell[     169] = 32'h0;  // 32'h9b9d7923;
    ram_cell[     170] = 32'h0;  // 32'h24d357c2;
    ram_cell[     171] = 32'h0;  // 32'h0457f6b0;
    ram_cell[     172] = 32'h0;  // 32'hc5a6a581;
    ram_cell[     173] = 32'h0;  // 32'h98cd8e1e;
    ram_cell[     174] = 32'h0;  // 32'h525b3917;
    ram_cell[     175] = 32'h0;  // 32'h283d2815;
    ram_cell[     176] = 32'h0;  // 32'h4c8cc969;
    ram_cell[     177] = 32'h0;  // 32'h04a344ed;
    ram_cell[     178] = 32'h0;  // 32'h0b40e089;
    ram_cell[     179] = 32'h0;  // 32'h0352d445;
    ram_cell[     180] = 32'h0;  // 32'h31898045;
    ram_cell[     181] = 32'h0;  // 32'h08b1f1ae;
    ram_cell[     182] = 32'h0;  // 32'h8ab00e06;
    ram_cell[     183] = 32'h0;  // 32'h5a82af0f;
    ram_cell[     184] = 32'h0;  // 32'h33e1fcc7;
    ram_cell[     185] = 32'h0;  // 32'hfcb56886;
    ram_cell[     186] = 32'h0;  // 32'h1018333e;
    ram_cell[     187] = 32'h0;  // 32'h3f2992a0;
    ram_cell[     188] = 32'h0;  // 32'h4eac07c6;
    ram_cell[     189] = 32'h0;  // 32'h84d51bc5;
    ram_cell[     190] = 32'h0;  // 32'h2f2ebaec;
    ram_cell[     191] = 32'h0;  // 32'hef1755c2;
    ram_cell[     192] = 32'h0;  // 32'hdd6f772e;
    ram_cell[     193] = 32'h0;  // 32'hc2780a53;
    ram_cell[     194] = 32'h0;  // 32'haa0eefca;
    ram_cell[     195] = 32'h0;  // 32'heeda0e76;
    ram_cell[     196] = 32'h0;  // 32'hd50b12b3;
    ram_cell[     197] = 32'h0;  // 32'h289257f0;
    ram_cell[     198] = 32'h0;  // 32'h3c2be22b;
    ram_cell[     199] = 32'h0;  // 32'hde22caf0;
    ram_cell[     200] = 32'h0;  // 32'haaacdea0;
    ram_cell[     201] = 32'h0;  // 32'hbffbe5d6;
    ram_cell[     202] = 32'h0;  // 32'hc403cd98;
    ram_cell[     203] = 32'h0;  // 32'h226bc821;
    ram_cell[     204] = 32'h0;  // 32'hdbf06b68;
    ram_cell[     205] = 32'h0;  // 32'h46c24393;
    ram_cell[     206] = 32'h0;  // 32'h2c0b8e95;
    ram_cell[     207] = 32'h0;  // 32'h1c8c88bf;
    ram_cell[     208] = 32'h0;  // 32'hb4b8a270;
    ram_cell[     209] = 32'h0;  // 32'h6f209db2;
    ram_cell[     210] = 32'h0;  // 32'h2404439a;
    ram_cell[     211] = 32'h0;  // 32'hda70c5d8;
    ram_cell[     212] = 32'h0;  // 32'h7918b178;
    ram_cell[     213] = 32'h0;  // 32'h75f686b9;
    ram_cell[     214] = 32'h0;  // 32'ha773c5de;
    ram_cell[     215] = 32'h0;  // 32'hdb4c3c36;
    ram_cell[     216] = 32'h0;  // 32'h35da439a;
    ram_cell[     217] = 32'h0;  // 32'hf8809f6f;
    ram_cell[     218] = 32'h0;  // 32'h8b7b8ec3;
    ram_cell[     219] = 32'h0;  // 32'hc69291f5;
    ram_cell[     220] = 32'h0;  // 32'h41156b9e;
    ram_cell[     221] = 32'h0;  // 32'h83620b9a;
    ram_cell[     222] = 32'h0;  // 32'hb26a533d;
    ram_cell[     223] = 32'h0;  // 32'h02784d72;
    ram_cell[     224] = 32'h0;  // 32'h71d7f509;
    ram_cell[     225] = 32'h0;  // 32'h720d6f6e;
    ram_cell[     226] = 32'h0;  // 32'hb95d00da;
    ram_cell[     227] = 32'h0;  // 32'hf27f249b;
    ram_cell[     228] = 32'h0;  // 32'he37928f0;
    ram_cell[     229] = 32'h0;  // 32'hce8a0804;
    ram_cell[     230] = 32'h0;  // 32'h4257bffb;
    ram_cell[     231] = 32'h0;  // 32'h152474f3;
    ram_cell[     232] = 32'h0;  // 32'h64976644;
    ram_cell[     233] = 32'h0;  // 32'hfb062104;
    ram_cell[     234] = 32'h0;  // 32'h13a84416;
    ram_cell[     235] = 32'h0;  // 32'h88b25276;
    ram_cell[     236] = 32'h0;  // 32'hdd3d552d;
    ram_cell[     237] = 32'h0;  // 32'h00368d43;
    ram_cell[     238] = 32'h0;  // 32'h80975443;
    ram_cell[     239] = 32'h0;  // 32'h8ecc0b1f;
    ram_cell[     240] = 32'h0;  // 32'h3eb857bb;
    ram_cell[     241] = 32'h0;  // 32'hd869bc59;
    ram_cell[     242] = 32'h0;  // 32'h9fa8ffcb;
    ram_cell[     243] = 32'h0;  // 32'h24faf85d;
    ram_cell[     244] = 32'h0;  // 32'hd1288628;
    ram_cell[     245] = 32'h0;  // 32'hbd0b075f;
    ram_cell[     246] = 32'h0;  // 32'hd23172f0;
    ram_cell[     247] = 32'h0;  // 32'h5ca55c0d;
    ram_cell[     248] = 32'h0;  // 32'h5c5a40f6;
    ram_cell[     249] = 32'h0;  // 32'h78d533e1;
    ram_cell[     250] = 32'h0;  // 32'h9594ecad;
    ram_cell[     251] = 32'h0;  // 32'h45ef7217;
    ram_cell[     252] = 32'h0;  // 32'hf3c66eeb;
    ram_cell[     253] = 32'h0;  // 32'h9b64259b;
    ram_cell[     254] = 32'h0;  // 32'h863f8358;
    ram_cell[     255] = 32'h0;  // 32'hecb3194b;
    // src matrix A
    ram_cell[     256] = 32'h2f22433c;
    ram_cell[     257] = 32'h93befdc8;
    ram_cell[     258] = 32'h2ef34452;
    ram_cell[     259] = 32'h65545b52;
    ram_cell[     260] = 32'hec02593b;
    ram_cell[     261] = 32'h8120ccf7;
    ram_cell[     262] = 32'h13eb59be;
    ram_cell[     263] = 32'h84b80941;
    ram_cell[     264] = 32'h8127597b;
    ram_cell[     265] = 32'h79f64b5f;
    ram_cell[     266] = 32'hf737368d;
    ram_cell[     267] = 32'h46b4a6c6;
    ram_cell[     268] = 32'h69152633;
    ram_cell[     269] = 32'h1dc0ab03;
    ram_cell[     270] = 32'h947715f7;
    ram_cell[     271] = 32'h6470ff4c;
    ram_cell[     272] = 32'hdbeb6e70;
    ram_cell[     273] = 32'h700c2edd;
    ram_cell[     274] = 32'hc31eab3a;
    ram_cell[     275] = 32'h7671a343;
    ram_cell[     276] = 32'h4fa96d20;
    ram_cell[     277] = 32'he774d470;
    ram_cell[     278] = 32'h8900f52e;
    ram_cell[     279] = 32'h0528ba1d;
    ram_cell[     280] = 32'h736c1351;
    ram_cell[     281] = 32'hd64d16a8;
    ram_cell[     282] = 32'h6d9f1c39;
    ram_cell[     283] = 32'hf585fe63;
    ram_cell[     284] = 32'h7b072b9a;
    ram_cell[     285] = 32'h55e10418;
    ram_cell[     286] = 32'h22e1cd04;
    ram_cell[     287] = 32'h6d22440a;
    ram_cell[     288] = 32'h719cdc62;
    ram_cell[     289] = 32'h1f0d7e44;
    ram_cell[     290] = 32'hccca1860;
    ram_cell[     291] = 32'h72e93bd2;
    ram_cell[     292] = 32'h827ebb2c;
    ram_cell[     293] = 32'h057b5306;
    ram_cell[     294] = 32'ha9cd9d49;
    ram_cell[     295] = 32'h196c9c4e;
    ram_cell[     296] = 32'h58988e87;
    ram_cell[     297] = 32'h32ea94c1;
    ram_cell[     298] = 32'h491e46d4;
    ram_cell[     299] = 32'hbfbaaa1f;
    ram_cell[     300] = 32'h10f70474;
    ram_cell[     301] = 32'hc6ad70c0;
    ram_cell[     302] = 32'hdfe83e12;
    ram_cell[     303] = 32'h0c353c1b;
    ram_cell[     304] = 32'h5f9c516b;
    ram_cell[     305] = 32'h79a15aa4;
    ram_cell[     306] = 32'he577874c;
    ram_cell[     307] = 32'h8833c850;
    ram_cell[     308] = 32'h674cb6d1;
    ram_cell[     309] = 32'h1458b613;
    ram_cell[     310] = 32'h340c18e0;
    ram_cell[     311] = 32'hd63a47dd;
    ram_cell[     312] = 32'hffcbeb3c;
    ram_cell[     313] = 32'h6652eef4;
    ram_cell[     314] = 32'h5d91686e;
    ram_cell[     315] = 32'he231ddaa;
    ram_cell[     316] = 32'h9e7b918e;
    ram_cell[     317] = 32'h34bfdb8d;
    ram_cell[     318] = 32'hdab521bd;
    ram_cell[     319] = 32'h8d90af0d;
    ram_cell[     320] = 32'h7bff4d54;
    ram_cell[     321] = 32'hfc5c44da;
    ram_cell[     322] = 32'hb078e70d;
    ram_cell[     323] = 32'hfc18c500;
    ram_cell[     324] = 32'h2cc6e66b;
    ram_cell[     325] = 32'h5b88b18d;
    ram_cell[     326] = 32'hf4d7debb;
    ram_cell[     327] = 32'hcc0babd2;
    ram_cell[     328] = 32'hbace89de;
    ram_cell[     329] = 32'h824b8bd3;
    ram_cell[     330] = 32'hc4d0a68c;
    ram_cell[     331] = 32'h64f3e55c;
    ram_cell[     332] = 32'h19f1a6d3;
    ram_cell[     333] = 32'hd2ccddf0;
    ram_cell[     334] = 32'ha9d29baa;
    ram_cell[     335] = 32'ha73e436d;
    ram_cell[     336] = 32'hcc2e2ca7;
    ram_cell[     337] = 32'h7f31909f;
    ram_cell[     338] = 32'hbc0521fb;
    ram_cell[     339] = 32'hd769d79a;
    ram_cell[     340] = 32'h64c44d09;
    ram_cell[     341] = 32'h0ea9479c;
    ram_cell[     342] = 32'hd0e2f1b2;
    ram_cell[     343] = 32'h7f242c29;
    ram_cell[     344] = 32'h7abe9388;
    ram_cell[     345] = 32'h22d57367;
    ram_cell[     346] = 32'h26cda775;
    ram_cell[     347] = 32'hd51a1c8f;
    ram_cell[     348] = 32'h86c8f0ba;
    ram_cell[     349] = 32'h0469d0db;
    ram_cell[     350] = 32'h3ec5d321;
    ram_cell[     351] = 32'hffe5cd44;
    ram_cell[     352] = 32'h380cf1d9;
    ram_cell[     353] = 32'h3c13929e;
    ram_cell[     354] = 32'hb35c0190;
    ram_cell[     355] = 32'h032c98ac;
    ram_cell[     356] = 32'h97272f8a;
    ram_cell[     357] = 32'h0b157cc0;
    ram_cell[     358] = 32'h48711f47;
    ram_cell[     359] = 32'h312ecff0;
    ram_cell[     360] = 32'hf33f6fe9;
    ram_cell[     361] = 32'h6ee94030;
    ram_cell[     362] = 32'heb27d6bc;
    ram_cell[     363] = 32'ha5d0355b;
    ram_cell[     364] = 32'h49445a93;
    ram_cell[     365] = 32'hfdef0411;
    ram_cell[     366] = 32'h4c03e08f;
    ram_cell[     367] = 32'h9e41a4b2;
    ram_cell[     368] = 32'h0d895fd9;
    ram_cell[     369] = 32'hbeae6cb8;
    ram_cell[     370] = 32'h225c75da;
    ram_cell[     371] = 32'he102da55;
    ram_cell[     372] = 32'h0ce68397;
    ram_cell[     373] = 32'h31304164;
    ram_cell[     374] = 32'h85a62d92;
    ram_cell[     375] = 32'hd59cdda2;
    ram_cell[     376] = 32'h9ac21d70;
    ram_cell[     377] = 32'hbc6cf657;
    ram_cell[     378] = 32'h2edb291a;
    ram_cell[     379] = 32'h40cc242c;
    ram_cell[     380] = 32'hdd33436d;
    ram_cell[     381] = 32'h8a63d9e3;
    ram_cell[     382] = 32'h91309a7b;
    ram_cell[     383] = 32'h3b5a978c;
    ram_cell[     384] = 32'h027490d7;
    ram_cell[     385] = 32'hb1b3673c;
    ram_cell[     386] = 32'h71576e03;
    ram_cell[     387] = 32'hb8c53b15;
    ram_cell[     388] = 32'h452221dc;
    ram_cell[     389] = 32'h8b3b0eff;
    ram_cell[     390] = 32'h5ea52389;
    ram_cell[     391] = 32'h2293a567;
    ram_cell[     392] = 32'h4a6a9895;
    ram_cell[     393] = 32'h98082310;
    ram_cell[     394] = 32'h4d8352ef;
    ram_cell[     395] = 32'h27efbf6d;
    ram_cell[     396] = 32'h97ed7b34;
    ram_cell[     397] = 32'hc3312f4d;
    ram_cell[     398] = 32'h84812085;
    ram_cell[     399] = 32'h37a8f1cf;
    ram_cell[     400] = 32'h6f86003f;
    ram_cell[     401] = 32'h9e5eb4d2;
    ram_cell[     402] = 32'h06539cc9;
    ram_cell[     403] = 32'h5d212af0;
    ram_cell[     404] = 32'ha4e3196a;
    ram_cell[     405] = 32'hddcc97e5;
    ram_cell[     406] = 32'h173f62a8;
    ram_cell[     407] = 32'h68ccb4f5;
    ram_cell[     408] = 32'hbc2558e2;
    ram_cell[     409] = 32'h2d6db3cd;
    ram_cell[     410] = 32'h7e890418;
    ram_cell[     411] = 32'hf6cc5230;
    ram_cell[     412] = 32'h7d4619f9;
    ram_cell[     413] = 32'hb66af771;
    ram_cell[     414] = 32'h86bd78ce;
    ram_cell[     415] = 32'hb4a1de00;
    ram_cell[     416] = 32'h9fa7ccdf;
    ram_cell[     417] = 32'h66ee6834;
    ram_cell[     418] = 32'he36b26b8;
    ram_cell[     419] = 32'hfba4710a;
    ram_cell[     420] = 32'h982ab136;
    ram_cell[     421] = 32'hce01fc80;
    ram_cell[     422] = 32'h6e495ae5;
    ram_cell[     423] = 32'hd28f684b;
    ram_cell[     424] = 32'hd6bc7435;
    ram_cell[     425] = 32'h8627e4e8;
    ram_cell[     426] = 32'hed186ba3;
    ram_cell[     427] = 32'h1d7225e3;
    ram_cell[     428] = 32'h3b059ea4;
    ram_cell[     429] = 32'h6621892d;
    ram_cell[     430] = 32'ha21f9f84;
    ram_cell[     431] = 32'h93b47ce5;
    ram_cell[     432] = 32'h997e602f;
    ram_cell[     433] = 32'h453ef143;
    ram_cell[     434] = 32'heea8e322;
    ram_cell[     435] = 32'hac10ac58;
    ram_cell[     436] = 32'he97c3f74;
    ram_cell[     437] = 32'h27810273;
    ram_cell[     438] = 32'hae4492e1;
    ram_cell[     439] = 32'h5a6b4e99;
    ram_cell[     440] = 32'h01e6e09f;
    ram_cell[     441] = 32'hc803fe49;
    ram_cell[     442] = 32'hde668a57;
    ram_cell[     443] = 32'hd8294669;
    ram_cell[     444] = 32'h5d6a0ee5;
    ram_cell[     445] = 32'h9ceea2d1;
    ram_cell[     446] = 32'h866fc7bb;
    ram_cell[     447] = 32'h7d88ab4c;
    ram_cell[     448] = 32'he2d86f04;
    ram_cell[     449] = 32'h607e0bbf;
    ram_cell[     450] = 32'h56950d67;
    ram_cell[     451] = 32'hbe1720d0;
    ram_cell[     452] = 32'hb31406af;
    ram_cell[     453] = 32'h51f5a705;
    ram_cell[     454] = 32'h6bc45205;
    ram_cell[     455] = 32'h0a8d0fea;
    ram_cell[     456] = 32'h7dada158;
    ram_cell[     457] = 32'hff88e854;
    ram_cell[     458] = 32'hb26ee3d8;
    ram_cell[     459] = 32'h5d06d20d;
    ram_cell[     460] = 32'ha9cec833;
    ram_cell[     461] = 32'h9de83aef;
    ram_cell[     462] = 32'h97d5a8a7;
    ram_cell[     463] = 32'hccc4de35;
    ram_cell[     464] = 32'hc43abc9d;
    ram_cell[     465] = 32'h898a02a8;
    ram_cell[     466] = 32'h96543468;
    ram_cell[     467] = 32'h9a4d04bb;
    ram_cell[     468] = 32'h43cb724c;
    ram_cell[     469] = 32'h0a22c87e;
    ram_cell[     470] = 32'h5734e472;
    ram_cell[     471] = 32'hae6f63ae;
    ram_cell[     472] = 32'hd1667b6a;
    ram_cell[     473] = 32'he7967712;
    ram_cell[     474] = 32'hacdd1d6e;
    ram_cell[     475] = 32'h8a6b32fa;
    ram_cell[     476] = 32'hb7d6c063;
    ram_cell[     477] = 32'hc3e19eaa;
    ram_cell[     478] = 32'h32311315;
    ram_cell[     479] = 32'hdff6cb63;
    ram_cell[     480] = 32'h2933d0cd;
    ram_cell[     481] = 32'hc6d4b91a;
    ram_cell[     482] = 32'h38aa0fd1;
    ram_cell[     483] = 32'h1be7e666;
    ram_cell[     484] = 32'hd7825837;
    ram_cell[     485] = 32'h4e1856a7;
    ram_cell[     486] = 32'h660e7089;
    ram_cell[     487] = 32'h642b3ff4;
    ram_cell[     488] = 32'h258da375;
    ram_cell[     489] = 32'h34e707bd;
    ram_cell[     490] = 32'h1150b566;
    ram_cell[     491] = 32'h330592e4;
    ram_cell[     492] = 32'hf961ac62;
    ram_cell[     493] = 32'h6d724e08;
    ram_cell[     494] = 32'hf54a6e93;
    ram_cell[     495] = 32'h821005fc;
    ram_cell[     496] = 32'hf5a75493;
    ram_cell[     497] = 32'hc42ccf89;
    ram_cell[     498] = 32'h657e524e;
    ram_cell[     499] = 32'hf38c6f8d;
    ram_cell[     500] = 32'h7b4f5020;
    ram_cell[     501] = 32'h0f4b5024;
    ram_cell[     502] = 32'h40cbf8e1;
    ram_cell[     503] = 32'h1654ede5;
    ram_cell[     504] = 32'ha72baac9;
    ram_cell[     505] = 32'h563a3b34;
    ram_cell[     506] = 32'hd1483bd8;
    ram_cell[     507] = 32'h4d03ac06;
    ram_cell[     508] = 32'h1258ca48;
    ram_cell[     509] = 32'h9a33f2a6;
    ram_cell[     510] = 32'h7b30b00c;
    ram_cell[     511] = 32'he450cb79;
    // src matrix B
    ram_cell[     512] = 32'hb45acdcd;
    ram_cell[     513] = 32'h074b282e;
    ram_cell[     514] = 32'h9950c1fb;
    ram_cell[     515] = 32'h0bed914a;
    ram_cell[     516] = 32'h51c49bf6;
    ram_cell[     517] = 32'ha30b9846;
    ram_cell[     518] = 32'h6984801b;
    ram_cell[     519] = 32'h393f442e;
    ram_cell[     520] = 32'h492aeb87;
    ram_cell[     521] = 32'h90662e3f;
    ram_cell[     522] = 32'hefb06188;
    ram_cell[     523] = 32'h20c58233;
    ram_cell[     524] = 32'h91adaf8c;
    ram_cell[     525] = 32'h2db6205c;
    ram_cell[     526] = 32'hd7d5935e;
    ram_cell[     527] = 32'h425b9ce1;
    ram_cell[     528] = 32'h7b204fc6;
    ram_cell[     529] = 32'h7d5af3cc;
    ram_cell[     530] = 32'h2def33c4;
    ram_cell[     531] = 32'hc532c0f2;
    ram_cell[     532] = 32'hafe4b1aa;
    ram_cell[     533] = 32'hf5e47009;
    ram_cell[     534] = 32'ha8818ab1;
    ram_cell[     535] = 32'hc774c801;
    ram_cell[     536] = 32'h02a94293;
    ram_cell[     537] = 32'h539e1dc7;
    ram_cell[     538] = 32'hbd5c9c71;
    ram_cell[     539] = 32'hc3227007;
    ram_cell[     540] = 32'hb4adc17f;
    ram_cell[     541] = 32'h150dded9;
    ram_cell[     542] = 32'hb29fa124;
    ram_cell[     543] = 32'hb7e91573;
    ram_cell[     544] = 32'h84f4a27f;
    ram_cell[     545] = 32'h82f37a19;
    ram_cell[     546] = 32'h41bc877e;
    ram_cell[     547] = 32'h6bcfd437;
    ram_cell[     548] = 32'h9d86cced;
    ram_cell[     549] = 32'hfec913b6;
    ram_cell[     550] = 32'h49dd1ddc;
    ram_cell[     551] = 32'h487a9821;
    ram_cell[     552] = 32'h4c29ceed;
    ram_cell[     553] = 32'hf5e48d4a;
    ram_cell[     554] = 32'h3ee324ea;
    ram_cell[     555] = 32'h6426b765;
    ram_cell[     556] = 32'h0f609553;
    ram_cell[     557] = 32'h1ea99085;
    ram_cell[     558] = 32'h4c202263;
    ram_cell[     559] = 32'hd626bc6d;
    ram_cell[     560] = 32'he702343d;
    ram_cell[     561] = 32'he472203d;
    ram_cell[     562] = 32'h5f34349d;
    ram_cell[     563] = 32'h3925bdf6;
    ram_cell[     564] = 32'h347a4323;
    ram_cell[     565] = 32'h68b7bafb;
    ram_cell[     566] = 32'h1f810c89;
    ram_cell[     567] = 32'h936ce08e;
    ram_cell[     568] = 32'h834c3376;
    ram_cell[     569] = 32'h59ab02b6;
    ram_cell[     570] = 32'h352c271c;
    ram_cell[     571] = 32'h50133314;
    ram_cell[     572] = 32'h98349d4b;
    ram_cell[     573] = 32'h22023d76;
    ram_cell[     574] = 32'h892f842a;
    ram_cell[     575] = 32'h4c862aff;
    ram_cell[     576] = 32'h9ac035a3;
    ram_cell[     577] = 32'hd38efc57;
    ram_cell[     578] = 32'h3605718f;
    ram_cell[     579] = 32'h5b73ea35;
    ram_cell[     580] = 32'hce9bf18e;
    ram_cell[     581] = 32'h4733759d;
    ram_cell[     582] = 32'h10bfe74b;
    ram_cell[     583] = 32'h99d2b659;
    ram_cell[     584] = 32'h12c6924c;
    ram_cell[     585] = 32'he867b151;
    ram_cell[     586] = 32'h5729d002;
    ram_cell[     587] = 32'hbf5fddc8;
    ram_cell[     588] = 32'h62f2b759;
    ram_cell[     589] = 32'h291495be;
    ram_cell[     590] = 32'h38fac543;
    ram_cell[     591] = 32'hda64eb70;
    ram_cell[     592] = 32'h32df3b6d;
    ram_cell[     593] = 32'hc27ef61d;
    ram_cell[     594] = 32'ha41a1a20;
    ram_cell[     595] = 32'hbddbfd0f;
    ram_cell[     596] = 32'h48db8e8b;
    ram_cell[     597] = 32'hb1e9381a;
    ram_cell[     598] = 32'hb8165152;
    ram_cell[     599] = 32'h9850257d;
    ram_cell[     600] = 32'he6e643c1;
    ram_cell[     601] = 32'h13492757;
    ram_cell[     602] = 32'h338218cb;
    ram_cell[     603] = 32'hf87f52c3;
    ram_cell[     604] = 32'hde9f6344;
    ram_cell[     605] = 32'h26351e56;
    ram_cell[     606] = 32'he59ae7fc;
    ram_cell[     607] = 32'hce7f3780;
    ram_cell[     608] = 32'h039acf12;
    ram_cell[     609] = 32'h6dca0231;
    ram_cell[     610] = 32'h2e53ae98;
    ram_cell[     611] = 32'h1c60901a;
    ram_cell[     612] = 32'h0744cbc3;
    ram_cell[     613] = 32'h85b7ad5c;
    ram_cell[     614] = 32'hdeacc350;
    ram_cell[     615] = 32'h36257b91;
    ram_cell[     616] = 32'hf3331a47;
    ram_cell[     617] = 32'h7f0a90d9;
    ram_cell[     618] = 32'h3e8155a2;
    ram_cell[     619] = 32'h249cd248;
    ram_cell[     620] = 32'hb5278579;
    ram_cell[     621] = 32'h0372d1ae;
    ram_cell[     622] = 32'he42eac23;
    ram_cell[     623] = 32'hf09e96b1;
    ram_cell[     624] = 32'h1d670014;
    ram_cell[     625] = 32'hf608a57a;
    ram_cell[     626] = 32'hfba0ad01;
    ram_cell[     627] = 32'h993d1b4f;
    ram_cell[     628] = 32'h791b9344;
    ram_cell[     629] = 32'hdf4f934f;
    ram_cell[     630] = 32'hb9b8e3be;
    ram_cell[     631] = 32'hc32a61d0;
    ram_cell[     632] = 32'h88d2782e;
    ram_cell[     633] = 32'hf7dcbb9d;
    ram_cell[     634] = 32'h6a986484;
    ram_cell[     635] = 32'hdceafa3a;
    ram_cell[     636] = 32'h5ddf5bd0;
    ram_cell[     637] = 32'hefcdce2c;
    ram_cell[     638] = 32'hd6eb33e1;
    ram_cell[     639] = 32'h7922cf74;
    ram_cell[     640] = 32'hfe7b21a8;
    ram_cell[     641] = 32'h5742be54;
    ram_cell[     642] = 32'h4d0ac54d;
    ram_cell[     643] = 32'ha83632b1;
    ram_cell[     644] = 32'h69c5d987;
    ram_cell[     645] = 32'h5d75a639;
    ram_cell[     646] = 32'ha5a44650;
    ram_cell[     647] = 32'h537da70f;
    ram_cell[     648] = 32'hb6f9d44a;
    ram_cell[     649] = 32'h8b97c0d9;
    ram_cell[     650] = 32'h54d55f24;
    ram_cell[     651] = 32'hb046a21f;
    ram_cell[     652] = 32'hc202aa86;
    ram_cell[     653] = 32'hbaa95d2a;
    ram_cell[     654] = 32'hf5de4176;
    ram_cell[     655] = 32'ha634e311;
    ram_cell[     656] = 32'hde80da27;
    ram_cell[     657] = 32'hb54905c5;
    ram_cell[     658] = 32'h5a300999;
    ram_cell[     659] = 32'ha2aac2ba;
    ram_cell[     660] = 32'h866ed42d;
    ram_cell[     661] = 32'h22424781;
    ram_cell[     662] = 32'h2883f35f;
    ram_cell[     663] = 32'h2f248f68;
    ram_cell[     664] = 32'h5feaf99e;
    ram_cell[     665] = 32'hb344d317;
    ram_cell[     666] = 32'h82179c9b;
    ram_cell[     667] = 32'h5499ce1e;
    ram_cell[     668] = 32'h06129e45;
    ram_cell[     669] = 32'ha8bfe470;
    ram_cell[     670] = 32'h4e933ef2;
    ram_cell[     671] = 32'he79c6208;
    ram_cell[     672] = 32'h9d28990c;
    ram_cell[     673] = 32'h65615728;
    ram_cell[     674] = 32'hededcd95;
    ram_cell[     675] = 32'hc2af8b54;
    ram_cell[     676] = 32'hc60f33f0;
    ram_cell[     677] = 32'h867d41f1;
    ram_cell[     678] = 32'hc54e5b2f;
    ram_cell[     679] = 32'h246a1714;
    ram_cell[     680] = 32'h3ba56110;
    ram_cell[     681] = 32'h9d4b42a5;
    ram_cell[     682] = 32'hce19bd1b;
    ram_cell[     683] = 32'h18d60c42;
    ram_cell[     684] = 32'hf7a10c1f;
    ram_cell[     685] = 32'hbe57af83;
    ram_cell[     686] = 32'h379a5cf6;
    ram_cell[     687] = 32'h528e99fc;
    ram_cell[     688] = 32'h2cd002a5;
    ram_cell[     689] = 32'he96111cd;
    ram_cell[     690] = 32'hb96dd399;
    ram_cell[     691] = 32'h4529e1bd;
    ram_cell[     692] = 32'h3c35b5ad;
    ram_cell[     693] = 32'h71677a6e;
    ram_cell[     694] = 32'h179d0f0b;
    ram_cell[     695] = 32'h2bb2df2f;
    ram_cell[     696] = 32'hae35f7fe;
    ram_cell[     697] = 32'hd5e92422;
    ram_cell[     698] = 32'hc91c34dd;
    ram_cell[     699] = 32'h423a3810;
    ram_cell[     700] = 32'h618a929f;
    ram_cell[     701] = 32'h77a01d67;
    ram_cell[     702] = 32'h705fee61;
    ram_cell[     703] = 32'he22c84cb;
    ram_cell[     704] = 32'h36738035;
    ram_cell[     705] = 32'hecb9e23b;
    ram_cell[     706] = 32'h6d80744b;
    ram_cell[     707] = 32'h1dcf1da0;
    ram_cell[     708] = 32'h84103eb1;
    ram_cell[     709] = 32'hc2a2498a;
    ram_cell[     710] = 32'h277cdbd9;
    ram_cell[     711] = 32'h3238896a;
    ram_cell[     712] = 32'h6abed080;
    ram_cell[     713] = 32'h8cdd8192;
    ram_cell[     714] = 32'h69c735e9;
    ram_cell[     715] = 32'hd8a636aa;
    ram_cell[     716] = 32'h44d1b76e;
    ram_cell[     717] = 32'h29ef36ae;
    ram_cell[     718] = 32'h8cdf5de7;
    ram_cell[     719] = 32'he931fc0f;
    ram_cell[     720] = 32'hd1f67112;
    ram_cell[     721] = 32'hb79389a9;
    ram_cell[     722] = 32'h791badaa;
    ram_cell[     723] = 32'hf7ecc9fa;
    ram_cell[     724] = 32'hc6ab7e26;
    ram_cell[     725] = 32'h5e6f8618;
    ram_cell[     726] = 32'hab1c3184;
    ram_cell[     727] = 32'h4c64d1c2;
    ram_cell[     728] = 32'h2ff491e7;
    ram_cell[     729] = 32'h056248b6;
    ram_cell[     730] = 32'hcaa4c752;
    ram_cell[     731] = 32'h7e4222aa;
    ram_cell[     732] = 32'h011b0b54;
    ram_cell[     733] = 32'h09841730;
    ram_cell[     734] = 32'h2ab9067e;
    ram_cell[     735] = 32'h6744d7e1;
    ram_cell[     736] = 32'h1690ba24;
    ram_cell[     737] = 32'hefc24b8d;
    ram_cell[     738] = 32'h5491e44a;
    ram_cell[     739] = 32'h4ab0a8b9;
    ram_cell[     740] = 32'h2e96a9c7;
    ram_cell[     741] = 32'hb76d535b;
    ram_cell[     742] = 32'hdbde8c9a;
    ram_cell[     743] = 32'h477b9532;
    ram_cell[     744] = 32'h112032ac;
    ram_cell[     745] = 32'h80465b6a;
    ram_cell[     746] = 32'h0453afb6;
    ram_cell[     747] = 32'h2ea360a6;
    ram_cell[     748] = 32'h4de16a15;
    ram_cell[     749] = 32'h16c96494;
    ram_cell[     750] = 32'hd1749d18;
    ram_cell[     751] = 32'h4ca81e49;
    ram_cell[     752] = 32'hf7a2f15f;
    ram_cell[     753] = 32'h61d94033;
    ram_cell[     754] = 32'hbf4a4f63;
    ram_cell[     755] = 32'hd83468bb;
    ram_cell[     756] = 32'hd57d4e1b;
    ram_cell[     757] = 32'h305568d1;
    ram_cell[     758] = 32'hf962f6f5;
    ram_cell[     759] = 32'h09f9c090;
    ram_cell[     760] = 32'hcd6c999f;
    ram_cell[     761] = 32'hd4064aae;
    ram_cell[     762] = 32'he7f126bc;
    ram_cell[     763] = 32'hc0eb8356;
    ram_cell[     764] = 32'he35f9502;
    ram_cell[     765] = 32'h9d1ec9a8;
    ram_cell[     766] = 32'h420adcaa;
    ram_cell[     767] = 32'h2f5e1ec0;
end

endmodule

