
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h0ee91e29;
    ram_cell[       1] = 32'h0;  // 32'hf6abc55b;
    ram_cell[       2] = 32'h0;  // 32'hd9af60f6;
    ram_cell[       3] = 32'h0;  // 32'hedad42a5;
    ram_cell[       4] = 32'h0;  // 32'hbec0d7f0;
    ram_cell[       5] = 32'h0;  // 32'h0bf06f68;
    ram_cell[       6] = 32'h0;  // 32'h45f2cdb8;
    ram_cell[       7] = 32'h0;  // 32'h09d2f0e8;
    ram_cell[       8] = 32'h0;  // 32'h45dcf81f;
    ram_cell[       9] = 32'h0;  // 32'h52644e6e;
    ram_cell[      10] = 32'h0;  // 32'hb57bb96f;
    ram_cell[      11] = 32'h0;  // 32'h624a521a;
    ram_cell[      12] = 32'h0;  // 32'h7ea45cd1;
    ram_cell[      13] = 32'h0;  // 32'h898c7b85;
    ram_cell[      14] = 32'h0;  // 32'hbb4f8a6f;
    ram_cell[      15] = 32'h0;  // 32'h23288065;
    ram_cell[      16] = 32'h0;  // 32'hc07ddb68;
    ram_cell[      17] = 32'h0;  // 32'h4ceccdca;
    ram_cell[      18] = 32'h0;  // 32'h11843cf2;
    ram_cell[      19] = 32'h0;  // 32'h6fb7fede;
    ram_cell[      20] = 32'h0;  // 32'ha604597c;
    ram_cell[      21] = 32'h0;  // 32'h6e124638;
    ram_cell[      22] = 32'h0;  // 32'he37ff407;
    ram_cell[      23] = 32'h0;  // 32'hc0edf216;
    ram_cell[      24] = 32'h0;  // 32'h85b83d28;
    ram_cell[      25] = 32'h0;  // 32'ha076d504;
    ram_cell[      26] = 32'h0;  // 32'he1a225da;
    ram_cell[      27] = 32'h0;  // 32'ha156a68b;
    ram_cell[      28] = 32'h0;  // 32'hc321bfac;
    ram_cell[      29] = 32'h0;  // 32'h38a66a86;
    ram_cell[      30] = 32'h0;  // 32'ha7e0feb5;
    ram_cell[      31] = 32'h0;  // 32'h46f8cec2;
    ram_cell[      32] = 32'h0;  // 32'h478d366e;
    ram_cell[      33] = 32'h0;  // 32'h0edd6f2c;
    ram_cell[      34] = 32'h0;  // 32'h9bd5e1c8;
    ram_cell[      35] = 32'h0;  // 32'hbe037cdc;
    ram_cell[      36] = 32'h0;  // 32'h365834c7;
    ram_cell[      37] = 32'h0;  // 32'h7b552514;
    ram_cell[      38] = 32'h0;  // 32'h53f51f3d;
    ram_cell[      39] = 32'h0;  // 32'hc1a11480;
    ram_cell[      40] = 32'h0;  // 32'hf2edbee2;
    ram_cell[      41] = 32'h0;  // 32'hc462e34c;
    ram_cell[      42] = 32'h0;  // 32'hd9ed6dbb;
    ram_cell[      43] = 32'h0;  // 32'h33456502;
    ram_cell[      44] = 32'h0;  // 32'h7cb8a692;
    ram_cell[      45] = 32'h0;  // 32'hea2e3a83;
    ram_cell[      46] = 32'h0;  // 32'h27e8c7b3;
    ram_cell[      47] = 32'h0;  // 32'h49fe7316;
    ram_cell[      48] = 32'h0;  // 32'h5bbbcb62;
    ram_cell[      49] = 32'h0;  // 32'h4d8fb720;
    ram_cell[      50] = 32'h0;  // 32'h0a5cf313;
    ram_cell[      51] = 32'h0;  // 32'h7a9d550a;
    ram_cell[      52] = 32'h0;  // 32'h1d90adee;
    ram_cell[      53] = 32'h0;  // 32'hf8fb61d9;
    ram_cell[      54] = 32'h0;  // 32'h95f71230;
    ram_cell[      55] = 32'h0;  // 32'hb83f8916;
    ram_cell[      56] = 32'h0;  // 32'h30c842fa;
    ram_cell[      57] = 32'h0;  // 32'h82b59a5b;
    ram_cell[      58] = 32'h0;  // 32'hc14f730a;
    ram_cell[      59] = 32'h0;  // 32'h59bf51ca;
    ram_cell[      60] = 32'h0;  // 32'hd27c71d1;
    ram_cell[      61] = 32'h0;  // 32'hc868517e;
    ram_cell[      62] = 32'h0;  // 32'h05223a54;
    ram_cell[      63] = 32'h0;  // 32'h795e9554;
    ram_cell[      64] = 32'h0;  // 32'h72c412aa;
    ram_cell[      65] = 32'h0;  // 32'h0c514a87;
    ram_cell[      66] = 32'h0;  // 32'h5a636e9b;
    ram_cell[      67] = 32'h0;  // 32'h25552468;
    ram_cell[      68] = 32'h0;  // 32'h6a3b4e6d;
    ram_cell[      69] = 32'h0;  // 32'h180382cf;
    ram_cell[      70] = 32'h0;  // 32'h5378ec0c;
    ram_cell[      71] = 32'h0;  // 32'h5d4aeb57;
    ram_cell[      72] = 32'h0;  // 32'h6f45f964;
    ram_cell[      73] = 32'h0;  // 32'h6383b1f6;
    ram_cell[      74] = 32'h0;  // 32'hd88ec217;
    ram_cell[      75] = 32'h0;  // 32'h4c8cacf2;
    ram_cell[      76] = 32'h0;  // 32'h76f3f0cb;
    ram_cell[      77] = 32'h0;  // 32'hba5cb555;
    ram_cell[      78] = 32'h0;  // 32'h41a7cb8a;
    ram_cell[      79] = 32'h0;  // 32'h7169ce13;
    ram_cell[      80] = 32'h0;  // 32'h6b4f5e49;
    ram_cell[      81] = 32'h0;  // 32'h13ad71ac;
    ram_cell[      82] = 32'h0;  // 32'he104e32c;
    ram_cell[      83] = 32'h0;  // 32'h8b9bdbad;
    ram_cell[      84] = 32'h0;  // 32'he67dd565;
    ram_cell[      85] = 32'h0;  // 32'h5d39ba5e;
    ram_cell[      86] = 32'h0;  // 32'h96714054;
    ram_cell[      87] = 32'h0;  // 32'h76c4c2fa;
    ram_cell[      88] = 32'h0;  // 32'h09e5e488;
    ram_cell[      89] = 32'h0;  // 32'hd1edb8a7;
    ram_cell[      90] = 32'h0;  // 32'h46aded7e;
    ram_cell[      91] = 32'h0;  // 32'h8a58cfe5;
    ram_cell[      92] = 32'h0;  // 32'h4fe418b9;
    ram_cell[      93] = 32'h0;  // 32'h154f6d69;
    ram_cell[      94] = 32'h0;  // 32'hae250bb6;
    ram_cell[      95] = 32'h0;  // 32'h8cf0949b;
    ram_cell[      96] = 32'h0;  // 32'h3cb0b125;
    ram_cell[      97] = 32'h0;  // 32'hbb146d4a;
    ram_cell[      98] = 32'h0;  // 32'hb31e2a11;
    ram_cell[      99] = 32'h0;  // 32'hf7e8260b;
    ram_cell[     100] = 32'h0;  // 32'hbcee7d67;
    ram_cell[     101] = 32'h0;  // 32'he3c1ad8b;
    ram_cell[     102] = 32'h0;  // 32'h807e7571;
    ram_cell[     103] = 32'h0;  // 32'h8180e29c;
    ram_cell[     104] = 32'h0;  // 32'h0b3ba778;
    ram_cell[     105] = 32'h0;  // 32'h216c71fb;
    ram_cell[     106] = 32'h0;  // 32'hd48854ed;
    ram_cell[     107] = 32'h0;  // 32'h07102568;
    ram_cell[     108] = 32'h0;  // 32'h1ff1dc44;
    ram_cell[     109] = 32'h0;  // 32'h924c6e27;
    ram_cell[     110] = 32'h0;  // 32'hb1be7e6f;
    ram_cell[     111] = 32'h0;  // 32'h807c4fa4;
    ram_cell[     112] = 32'h0;  // 32'h43d436cd;
    ram_cell[     113] = 32'h0;  // 32'h3d68ebd2;
    ram_cell[     114] = 32'h0;  // 32'ha88981fe;
    ram_cell[     115] = 32'h0;  // 32'hfc1ffb2d;
    ram_cell[     116] = 32'h0;  // 32'h184df444;
    ram_cell[     117] = 32'h0;  // 32'h40eabea0;
    ram_cell[     118] = 32'h0;  // 32'hdde725e4;
    ram_cell[     119] = 32'h0;  // 32'h4e76624f;
    ram_cell[     120] = 32'h0;  // 32'h79d2acbd;
    ram_cell[     121] = 32'h0;  // 32'hee9719fd;
    ram_cell[     122] = 32'h0;  // 32'h9cdddc46;
    ram_cell[     123] = 32'h0;  // 32'h479df452;
    ram_cell[     124] = 32'h0;  // 32'hc9d3302c;
    ram_cell[     125] = 32'h0;  // 32'h55ff1f8c;
    ram_cell[     126] = 32'h0;  // 32'he9d8820f;
    ram_cell[     127] = 32'h0;  // 32'h1a7786fc;
    ram_cell[     128] = 32'h0;  // 32'h15392fc4;
    ram_cell[     129] = 32'h0;  // 32'h4b54da2f;
    ram_cell[     130] = 32'h0;  // 32'h68da69b3;
    ram_cell[     131] = 32'h0;  // 32'ha012e3e5;
    ram_cell[     132] = 32'h0;  // 32'h85af6d6c;
    ram_cell[     133] = 32'h0;  // 32'h5937b43b;
    ram_cell[     134] = 32'h0;  // 32'hd98e1ebe;
    ram_cell[     135] = 32'h0;  // 32'h50cbdb27;
    ram_cell[     136] = 32'h0;  // 32'h491d3453;
    ram_cell[     137] = 32'h0;  // 32'hc7767e46;
    ram_cell[     138] = 32'h0;  // 32'hfe584e60;
    ram_cell[     139] = 32'h0;  // 32'h5068b01b;
    ram_cell[     140] = 32'h0;  // 32'h4b7ffe28;
    ram_cell[     141] = 32'h0;  // 32'h722d0cff;
    ram_cell[     142] = 32'h0;  // 32'h089b160b;
    ram_cell[     143] = 32'h0;  // 32'he4afa66c;
    ram_cell[     144] = 32'h0;  // 32'h96dfac2a;
    ram_cell[     145] = 32'h0;  // 32'h7641d47d;
    ram_cell[     146] = 32'h0;  // 32'hc500d2ab;
    ram_cell[     147] = 32'h0;  // 32'h81af69b2;
    ram_cell[     148] = 32'h0;  // 32'hd6b3ce26;
    ram_cell[     149] = 32'h0;  // 32'h96284645;
    ram_cell[     150] = 32'h0;  // 32'h873424c8;
    ram_cell[     151] = 32'h0;  // 32'h5e7852a1;
    ram_cell[     152] = 32'h0;  // 32'h67bc575e;
    ram_cell[     153] = 32'h0;  // 32'he7d71e84;
    ram_cell[     154] = 32'h0;  // 32'h395056c5;
    ram_cell[     155] = 32'h0;  // 32'h3bcd09b3;
    ram_cell[     156] = 32'h0;  // 32'h656ae2fe;
    ram_cell[     157] = 32'h0;  // 32'h9a8af298;
    ram_cell[     158] = 32'h0;  // 32'hf43c5b69;
    ram_cell[     159] = 32'h0;  // 32'hc227ede2;
    ram_cell[     160] = 32'h0;  // 32'h7c96a833;
    ram_cell[     161] = 32'h0;  // 32'hc45bc461;
    ram_cell[     162] = 32'h0;  // 32'hd9ef5711;
    ram_cell[     163] = 32'h0;  // 32'h8c5a1ee6;
    ram_cell[     164] = 32'h0;  // 32'h62140631;
    ram_cell[     165] = 32'h0;  // 32'h0cd62988;
    ram_cell[     166] = 32'h0;  // 32'hed1ad81a;
    ram_cell[     167] = 32'h0;  // 32'h54eacbf8;
    ram_cell[     168] = 32'h0;  // 32'h94c8509b;
    ram_cell[     169] = 32'h0;  // 32'h5693006b;
    ram_cell[     170] = 32'h0;  // 32'hd56bdfe0;
    ram_cell[     171] = 32'h0;  // 32'h937c4fce;
    ram_cell[     172] = 32'h0;  // 32'h1b32e39f;
    ram_cell[     173] = 32'h0;  // 32'h41b33ef3;
    ram_cell[     174] = 32'h0;  // 32'h03a83c84;
    ram_cell[     175] = 32'h0;  // 32'hea86875b;
    ram_cell[     176] = 32'h0;  // 32'h93ae224f;
    ram_cell[     177] = 32'h0;  // 32'hd01e2e54;
    ram_cell[     178] = 32'h0;  // 32'h2e9d1eac;
    ram_cell[     179] = 32'h0;  // 32'h659f7bf5;
    ram_cell[     180] = 32'h0;  // 32'h0a39a386;
    ram_cell[     181] = 32'h0;  // 32'h0220e0d7;
    ram_cell[     182] = 32'h0;  // 32'h604c5b2f;
    ram_cell[     183] = 32'h0;  // 32'hb782bfb2;
    ram_cell[     184] = 32'h0;  // 32'h6be562b7;
    ram_cell[     185] = 32'h0;  // 32'h32a42729;
    ram_cell[     186] = 32'h0;  // 32'h5d862ad8;
    ram_cell[     187] = 32'h0;  // 32'h8fef4b2e;
    ram_cell[     188] = 32'h0;  // 32'h611b458d;
    ram_cell[     189] = 32'h0;  // 32'hcd435ed7;
    ram_cell[     190] = 32'h0;  // 32'h32cb9075;
    ram_cell[     191] = 32'h0;  // 32'h7d281891;
    ram_cell[     192] = 32'h0;  // 32'hcfa64c39;
    ram_cell[     193] = 32'h0;  // 32'h1fc77f0b;
    ram_cell[     194] = 32'h0;  // 32'hd07a8cc0;
    ram_cell[     195] = 32'h0;  // 32'h29018919;
    ram_cell[     196] = 32'h0;  // 32'h2c29ef87;
    ram_cell[     197] = 32'h0;  // 32'hd4434da6;
    ram_cell[     198] = 32'h0;  // 32'h6969dd97;
    ram_cell[     199] = 32'h0;  // 32'h26a8f4ca;
    ram_cell[     200] = 32'h0;  // 32'ha38da532;
    ram_cell[     201] = 32'h0;  // 32'h6590e8e8;
    ram_cell[     202] = 32'h0;  // 32'h61e49313;
    ram_cell[     203] = 32'h0;  // 32'h0422ddc3;
    ram_cell[     204] = 32'h0;  // 32'ha4da3743;
    ram_cell[     205] = 32'h0;  // 32'h89bcecb5;
    ram_cell[     206] = 32'h0;  // 32'h544ae086;
    ram_cell[     207] = 32'h0;  // 32'hd6794d29;
    ram_cell[     208] = 32'h0;  // 32'h712b3156;
    ram_cell[     209] = 32'h0;  // 32'h80db0d3e;
    ram_cell[     210] = 32'h0;  // 32'h354cdfac;
    ram_cell[     211] = 32'h0;  // 32'h6d88168a;
    ram_cell[     212] = 32'h0;  // 32'h557070ca;
    ram_cell[     213] = 32'h0;  // 32'hccc507ab;
    ram_cell[     214] = 32'h0;  // 32'hebaf9d3b;
    ram_cell[     215] = 32'h0;  // 32'h05b2c165;
    ram_cell[     216] = 32'h0;  // 32'hb7097cdc;
    ram_cell[     217] = 32'h0;  // 32'h6973a698;
    ram_cell[     218] = 32'h0;  // 32'h73c3789c;
    ram_cell[     219] = 32'h0;  // 32'h5b0092bc;
    ram_cell[     220] = 32'h0;  // 32'h34b3f8b4;
    ram_cell[     221] = 32'h0;  // 32'h6befe236;
    ram_cell[     222] = 32'h0;  // 32'h103bf5a5;
    ram_cell[     223] = 32'h0;  // 32'h33db3a13;
    ram_cell[     224] = 32'h0;  // 32'h24c734c6;
    ram_cell[     225] = 32'h0;  // 32'h2d77f8b6;
    ram_cell[     226] = 32'h0;  // 32'hf5414ea3;
    ram_cell[     227] = 32'h0;  // 32'hd828759a;
    ram_cell[     228] = 32'h0;  // 32'ha06b061c;
    ram_cell[     229] = 32'h0;  // 32'hbc4184cc;
    ram_cell[     230] = 32'h0;  // 32'h93a26fb5;
    ram_cell[     231] = 32'h0;  // 32'h368546bb;
    ram_cell[     232] = 32'h0;  // 32'h4060f4ef;
    ram_cell[     233] = 32'h0;  // 32'hfdc78bd4;
    ram_cell[     234] = 32'h0;  // 32'h700d69b6;
    ram_cell[     235] = 32'h0;  // 32'hf0bc72bc;
    ram_cell[     236] = 32'h0;  // 32'hf7afa0a5;
    ram_cell[     237] = 32'h0;  // 32'h3c3c4c0c;
    ram_cell[     238] = 32'h0;  // 32'hdd24138f;
    ram_cell[     239] = 32'h0;  // 32'h30efebf7;
    ram_cell[     240] = 32'h0;  // 32'hd377dbc0;
    ram_cell[     241] = 32'h0;  // 32'hde1c377d;
    ram_cell[     242] = 32'h0;  // 32'h07282509;
    ram_cell[     243] = 32'h0;  // 32'heedf87b4;
    ram_cell[     244] = 32'h0;  // 32'h5b729e41;
    ram_cell[     245] = 32'h0;  // 32'h22b7b089;
    ram_cell[     246] = 32'h0;  // 32'h2211d512;
    ram_cell[     247] = 32'h0;  // 32'ha4ff778e;
    ram_cell[     248] = 32'h0;  // 32'hdd0e3f37;
    ram_cell[     249] = 32'h0;  // 32'h61f54fce;
    ram_cell[     250] = 32'h0;  // 32'haf9164e0;
    ram_cell[     251] = 32'h0;  // 32'h8e85c231;
    ram_cell[     252] = 32'h0;  // 32'hcd7dc990;
    ram_cell[     253] = 32'h0;  // 32'hd351ab60;
    ram_cell[     254] = 32'h0;  // 32'h79f41d8e;
    ram_cell[     255] = 32'h0;  // 32'hfe289977;
    // src matrix A
    ram_cell[     256] = 32'h69efb9a9;
    ram_cell[     257] = 32'h4db1c6ab;
    ram_cell[     258] = 32'h72edf36e;
    ram_cell[     259] = 32'hc3d40dcd;
    ram_cell[     260] = 32'h3825b927;
    ram_cell[     261] = 32'hd7cbe275;
    ram_cell[     262] = 32'ha599a069;
    ram_cell[     263] = 32'hce024147;
    ram_cell[     264] = 32'hba663fbb;
    ram_cell[     265] = 32'hde4bff19;
    ram_cell[     266] = 32'h7b292645;
    ram_cell[     267] = 32'h10a388d5;
    ram_cell[     268] = 32'h1059ca0d;
    ram_cell[     269] = 32'ha97c3029;
    ram_cell[     270] = 32'h6aab6d6d;
    ram_cell[     271] = 32'hfce841f3;
    ram_cell[     272] = 32'h1d3e759d;
    ram_cell[     273] = 32'he6ef94ee;
    ram_cell[     274] = 32'hfc2af7f0;
    ram_cell[     275] = 32'h5a84f6ad;
    ram_cell[     276] = 32'h9374f2f5;
    ram_cell[     277] = 32'h9716c7c4;
    ram_cell[     278] = 32'ha2086da5;
    ram_cell[     279] = 32'h5b83c50e;
    ram_cell[     280] = 32'hea4e6467;
    ram_cell[     281] = 32'h6fc6b8f7;
    ram_cell[     282] = 32'h672683df;
    ram_cell[     283] = 32'h8cd0f907;
    ram_cell[     284] = 32'h3e8d623a;
    ram_cell[     285] = 32'h9ccf28f8;
    ram_cell[     286] = 32'h043a6835;
    ram_cell[     287] = 32'h437202b6;
    ram_cell[     288] = 32'h50012fda;
    ram_cell[     289] = 32'h2d453733;
    ram_cell[     290] = 32'h16ca90df;
    ram_cell[     291] = 32'h1a497013;
    ram_cell[     292] = 32'hf889389f;
    ram_cell[     293] = 32'hb5e6022d;
    ram_cell[     294] = 32'he212a86e;
    ram_cell[     295] = 32'hd6a15bbf;
    ram_cell[     296] = 32'h57f5d893;
    ram_cell[     297] = 32'h4857b2e3;
    ram_cell[     298] = 32'hd45a36b0;
    ram_cell[     299] = 32'hf1ca2a8b;
    ram_cell[     300] = 32'h010ec5ee;
    ram_cell[     301] = 32'h0d07c41b;
    ram_cell[     302] = 32'he1099e76;
    ram_cell[     303] = 32'hff7d0baa;
    ram_cell[     304] = 32'h0199cfb7;
    ram_cell[     305] = 32'h7003ec67;
    ram_cell[     306] = 32'hb9414fda;
    ram_cell[     307] = 32'hfd3acf7e;
    ram_cell[     308] = 32'hf15d93c1;
    ram_cell[     309] = 32'h0a321e1d;
    ram_cell[     310] = 32'h2bc8a9ff;
    ram_cell[     311] = 32'h711975f2;
    ram_cell[     312] = 32'h1c20e397;
    ram_cell[     313] = 32'hd54f1cd8;
    ram_cell[     314] = 32'ha6fc776f;
    ram_cell[     315] = 32'he5bd0e4e;
    ram_cell[     316] = 32'hb2435638;
    ram_cell[     317] = 32'h595bb515;
    ram_cell[     318] = 32'h4a44715b;
    ram_cell[     319] = 32'h0285e73a;
    ram_cell[     320] = 32'h087b88c8;
    ram_cell[     321] = 32'hfceeb1e8;
    ram_cell[     322] = 32'he97e60ca;
    ram_cell[     323] = 32'h1e5326ac;
    ram_cell[     324] = 32'h5e604e04;
    ram_cell[     325] = 32'hff8792bf;
    ram_cell[     326] = 32'h4fc0c50f;
    ram_cell[     327] = 32'he49c441e;
    ram_cell[     328] = 32'h3d91a332;
    ram_cell[     329] = 32'h2f0af157;
    ram_cell[     330] = 32'h67d94f06;
    ram_cell[     331] = 32'h8d37c77e;
    ram_cell[     332] = 32'h6f43e84d;
    ram_cell[     333] = 32'h4b0afa68;
    ram_cell[     334] = 32'hd4deff2f;
    ram_cell[     335] = 32'h050ce59a;
    ram_cell[     336] = 32'hcc6c473a;
    ram_cell[     337] = 32'h859fc93c;
    ram_cell[     338] = 32'h4161a65e;
    ram_cell[     339] = 32'hdc615f23;
    ram_cell[     340] = 32'h659319f8;
    ram_cell[     341] = 32'h18c2cbb7;
    ram_cell[     342] = 32'h2fd84cfd;
    ram_cell[     343] = 32'h360f7cee;
    ram_cell[     344] = 32'h263a2499;
    ram_cell[     345] = 32'ha1a67ef6;
    ram_cell[     346] = 32'h8639b4b6;
    ram_cell[     347] = 32'h1d14bd99;
    ram_cell[     348] = 32'haa2f880b;
    ram_cell[     349] = 32'h10633797;
    ram_cell[     350] = 32'h42cb1ecb;
    ram_cell[     351] = 32'h50368f17;
    ram_cell[     352] = 32'h8e5325d8;
    ram_cell[     353] = 32'h74db17fe;
    ram_cell[     354] = 32'hafcaeef4;
    ram_cell[     355] = 32'h056b82cc;
    ram_cell[     356] = 32'h5ffe7291;
    ram_cell[     357] = 32'h6dca9aba;
    ram_cell[     358] = 32'hee68ba7e;
    ram_cell[     359] = 32'he4ef96dc;
    ram_cell[     360] = 32'h754f7317;
    ram_cell[     361] = 32'hdfcbeac3;
    ram_cell[     362] = 32'had99bd8e;
    ram_cell[     363] = 32'h4e308f0c;
    ram_cell[     364] = 32'h80f7bd9b;
    ram_cell[     365] = 32'h82767d74;
    ram_cell[     366] = 32'h5111aa5f;
    ram_cell[     367] = 32'ha0aa5574;
    ram_cell[     368] = 32'h8a1fd1a6;
    ram_cell[     369] = 32'h28c24b3e;
    ram_cell[     370] = 32'ha1f54027;
    ram_cell[     371] = 32'h5a6e12d2;
    ram_cell[     372] = 32'hcf895520;
    ram_cell[     373] = 32'h8dfc44fe;
    ram_cell[     374] = 32'h1c776680;
    ram_cell[     375] = 32'h691b14bf;
    ram_cell[     376] = 32'h35bcd292;
    ram_cell[     377] = 32'hc3534087;
    ram_cell[     378] = 32'h2ef1e770;
    ram_cell[     379] = 32'h0c996a7b;
    ram_cell[     380] = 32'he40616e1;
    ram_cell[     381] = 32'h02fa02d8;
    ram_cell[     382] = 32'h0434f227;
    ram_cell[     383] = 32'h3ea74eed;
    ram_cell[     384] = 32'haeebb614;
    ram_cell[     385] = 32'h4cf6f208;
    ram_cell[     386] = 32'hafc73cb1;
    ram_cell[     387] = 32'h1c44b425;
    ram_cell[     388] = 32'h723c985f;
    ram_cell[     389] = 32'h80a780ab;
    ram_cell[     390] = 32'ha11d6f56;
    ram_cell[     391] = 32'hb6a166ef;
    ram_cell[     392] = 32'h4285cc28;
    ram_cell[     393] = 32'hf1166341;
    ram_cell[     394] = 32'he5158850;
    ram_cell[     395] = 32'h8ba66a35;
    ram_cell[     396] = 32'hee8460ea;
    ram_cell[     397] = 32'hca986295;
    ram_cell[     398] = 32'h184fb568;
    ram_cell[     399] = 32'haef6a73c;
    ram_cell[     400] = 32'h5fb18b74;
    ram_cell[     401] = 32'h010eb1e3;
    ram_cell[     402] = 32'h2f2bfdac;
    ram_cell[     403] = 32'h5e35f4a7;
    ram_cell[     404] = 32'hacf56a1b;
    ram_cell[     405] = 32'hc2069c64;
    ram_cell[     406] = 32'h2abb17a1;
    ram_cell[     407] = 32'h20edab94;
    ram_cell[     408] = 32'hb8ad50b2;
    ram_cell[     409] = 32'h196a6193;
    ram_cell[     410] = 32'hef564b83;
    ram_cell[     411] = 32'h4ecd4de9;
    ram_cell[     412] = 32'h7ff1e05f;
    ram_cell[     413] = 32'h9f227b91;
    ram_cell[     414] = 32'he0d11fb9;
    ram_cell[     415] = 32'ha06489d0;
    ram_cell[     416] = 32'hfbdbd13b;
    ram_cell[     417] = 32'h52e9a05a;
    ram_cell[     418] = 32'h49bc8a80;
    ram_cell[     419] = 32'h98e3b8fe;
    ram_cell[     420] = 32'h00614d64;
    ram_cell[     421] = 32'h1e4757f5;
    ram_cell[     422] = 32'h95beab2c;
    ram_cell[     423] = 32'h930a0314;
    ram_cell[     424] = 32'h58dc3cbf;
    ram_cell[     425] = 32'h28b2c17e;
    ram_cell[     426] = 32'h33467b9e;
    ram_cell[     427] = 32'hc62930af;
    ram_cell[     428] = 32'hb4867a92;
    ram_cell[     429] = 32'h23048d54;
    ram_cell[     430] = 32'h1f08d916;
    ram_cell[     431] = 32'h37b4add2;
    ram_cell[     432] = 32'h0d586fbb;
    ram_cell[     433] = 32'h1f5ef08f;
    ram_cell[     434] = 32'hd34e7961;
    ram_cell[     435] = 32'h7165895b;
    ram_cell[     436] = 32'hfe3c67b0;
    ram_cell[     437] = 32'hc4c73046;
    ram_cell[     438] = 32'hcc89c0c7;
    ram_cell[     439] = 32'h6c22b03d;
    ram_cell[     440] = 32'h425cf7be;
    ram_cell[     441] = 32'h0a0bbe1f;
    ram_cell[     442] = 32'he3c42ba6;
    ram_cell[     443] = 32'h352176fd;
    ram_cell[     444] = 32'hbfdc6c32;
    ram_cell[     445] = 32'h487b7ca9;
    ram_cell[     446] = 32'h70a3755d;
    ram_cell[     447] = 32'he34a8844;
    ram_cell[     448] = 32'h5d0047d2;
    ram_cell[     449] = 32'h5d90573c;
    ram_cell[     450] = 32'hf211a1f8;
    ram_cell[     451] = 32'h7a217121;
    ram_cell[     452] = 32'hec418c8c;
    ram_cell[     453] = 32'h8d54c148;
    ram_cell[     454] = 32'heb002965;
    ram_cell[     455] = 32'h950c8885;
    ram_cell[     456] = 32'h80f89a76;
    ram_cell[     457] = 32'hd134f6b7;
    ram_cell[     458] = 32'h1c5e884a;
    ram_cell[     459] = 32'h8dc2302a;
    ram_cell[     460] = 32'he49fb8d2;
    ram_cell[     461] = 32'h6152998c;
    ram_cell[     462] = 32'h57ea8765;
    ram_cell[     463] = 32'hd5746ee3;
    ram_cell[     464] = 32'hdb7b72ef;
    ram_cell[     465] = 32'h7a2dfcda;
    ram_cell[     466] = 32'h2ac865e0;
    ram_cell[     467] = 32'hef7363f1;
    ram_cell[     468] = 32'hbd01b254;
    ram_cell[     469] = 32'h23e119f2;
    ram_cell[     470] = 32'h89ddce24;
    ram_cell[     471] = 32'hb68876ce;
    ram_cell[     472] = 32'hdd178da1;
    ram_cell[     473] = 32'h2529ea1b;
    ram_cell[     474] = 32'h3a044edc;
    ram_cell[     475] = 32'h7bd8e605;
    ram_cell[     476] = 32'h09be791a;
    ram_cell[     477] = 32'h70eb9534;
    ram_cell[     478] = 32'hfe3f4f95;
    ram_cell[     479] = 32'h77e19ccf;
    ram_cell[     480] = 32'h8866d524;
    ram_cell[     481] = 32'he0c8b6d5;
    ram_cell[     482] = 32'hd2616618;
    ram_cell[     483] = 32'hc28a1880;
    ram_cell[     484] = 32'h1e712a28;
    ram_cell[     485] = 32'h0cc8e139;
    ram_cell[     486] = 32'h7175bab1;
    ram_cell[     487] = 32'h608cf7d7;
    ram_cell[     488] = 32'h2c0fdcc7;
    ram_cell[     489] = 32'h70e5ece2;
    ram_cell[     490] = 32'h8ef9af06;
    ram_cell[     491] = 32'h6bcd8934;
    ram_cell[     492] = 32'h7cf4d550;
    ram_cell[     493] = 32'hde3cd397;
    ram_cell[     494] = 32'ha8d425b3;
    ram_cell[     495] = 32'hdf7c96f9;
    ram_cell[     496] = 32'h4316dad5;
    ram_cell[     497] = 32'h56691132;
    ram_cell[     498] = 32'h111df645;
    ram_cell[     499] = 32'h1b056ae7;
    ram_cell[     500] = 32'h25820daf;
    ram_cell[     501] = 32'ha875ad1b;
    ram_cell[     502] = 32'hc6e007b0;
    ram_cell[     503] = 32'h6832b8c8;
    ram_cell[     504] = 32'h627d3049;
    ram_cell[     505] = 32'h162b8151;
    ram_cell[     506] = 32'h03edc906;
    ram_cell[     507] = 32'h65985573;
    ram_cell[     508] = 32'hdfc868c8;
    ram_cell[     509] = 32'h0b25a41b;
    ram_cell[     510] = 32'h176b46fe;
    ram_cell[     511] = 32'h526d335e;
    // src matrix B
    ram_cell[     512] = 32'h6eed6478;
    ram_cell[     513] = 32'h8d1d2a45;
    ram_cell[     514] = 32'haca7bfd3;
    ram_cell[     515] = 32'h23d9a93b;
    ram_cell[     516] = 32'h72c58a96;
    ram_cell[     517] = 32'h8ec63441;
    ram_cell[     518] = 32'h145fd615;
    ram_cell[     519] = 32'h2425bb76;
    ram_cell[     520] = 32'h41e86019;
    ram_cell[     521] = 32'hbf94f718;
    ram_cell[     522] = 32'hf367f33b;
    ram_cell[     523] = 32'he5322031;
    ram_cell[     524] = 32'h4f1bf1da;
    ram_cell[     525] = 32'h40c978b4;
    ram_cell[     526] = 32'h1ae49796;
    ram_cell[     527] = 32'h5742bead;
    ram_cell[     528] = 32'h8fe458a4;
    ram_cell[     529] = 32'h3b968df1;
    ram_cell[     530] = 32'hf9f6d364;
    ram_cell[     531] = 32'h9c6b5988;
    ram_cell[     532] = 32'h42d848f7;
    ram_cell[     533] = 32'hb82c72b3;
    ram_cell[     534] = 32'h26d96a11;
    ram_cell[     535] = 32'hd1e82984;
    ram_cell[     536] = 32'h08c71007;
    ram_cell[     537] = 32'hadae488a;
    ram_cell[     538] = 32'ha96ab33e;
    ram_cell[     539] = 32'he8697712;
    ram_cell[     540] = 32'h385d08bd;
    ram_cell[     541] = 32'h4a6510ff;
    ram_cell[     542] = 32'hf84107e7;
    ram_cell[     543] = 32'h7f2623c2;
    ram_cell[     544] = 32'h1d28d763;
    ram_cell[     545] = 32'h302a5291;
    ram_cell[     546] = 32'h4f3a02a2;
    ram_cell[     547] = 32'he2b92e5c;
    ram_cell[     548] = 32'h0b4ae707;
    ram_cell[     549] = 32'h9f1d45d2;
    ram_cell[     550] = 32'h27fa24c3;
    ram_cell[     551] = 32'ha62cd5ba;
    ram_cell[     552] = 32'hd88e8c01;
    ram_cell[     553] = 32'h7eebe4b9;
    ram_cell[     554] = 32'hb497637e;
    ram_cell[     555] = 32'hd6623ce4;
    ram_cell[     556] = 32'h11138d6c;
    ram_cell[     557] = 32'hd8190b03;
    ram_cell[     558] = 32'hcdc83316;
    ram_cell[     559] = 32'h369c3d62;
    ram_cell[     560] = 32'h2afecfed;
    ram_cell[     561] = 32'hf94512ee;
    ram_cell[     562] = 32'hdf957be2;
    ram_cell[     563] = 32'h78ba8463;
    ram_cell[     564] = 32'h5af25872;
    ram_cell[     565] = 32'h542d79ff;
    ram_cell[     566] = 32'h0bf3f627;
    ram_cell[     567] = 32'h528652e0;
    ram_cell[     568] = 32'h574d3421;
    ram_cell[     569] = 32'h5ee9b6d5;
    ram_cell[     570] = 32'hac29b81d;
    ram_cell[     571] = 32'h63d1cb07;
    ram_cell[     572] = 32'h74e85db8;
    ram_cell[     573] = 32'hec69b4fe;
    ram_cell[     574] = 32'h57797879;
    ram_cell[     575] = 32'hac3d9d6e;
    ram_cell[     576] = 32'hb3dd4153;
    ram_cell[     577] = 32'he90bc822;
    ram_cell[     578] = 32'h2d421360;
    ram_cell[     579] = 32'h904aaef4;
    ram_cell[     580] = 32'h5335c541;
    ram_cell[     581] = 32'hb317f5e0;
    ram_cell[     582] = 32'hb1308c2c;
    ram_cell[     583] = 32'h3b107be3;
    ram_cell[     584] = 32'h029a3eee;
    ram_cell[     585] = 32'h9bed095e;
    ram_cell[     586] = 32'hd1b1bcde;
    ram_cell[     587] = 32'h49ae7cd2;
    ram_cell[     588] = 32'h49028fb1;
    ram_cell[     589] = 32'h269c77cd;
    ram_cell[     590] = 32'h8f5d4091;
    ram_cell[     591] = 32'h8443fe16;
    ram_cell[     592] = 32'h4e7b11c0;
    ram_cell[     593] = 32'h636fa109;
    ram_cell[     594] = 32'h0c128014;
    ram_cell[     595] = 32'h7feab45e;
    ram_cell[     596] = 32'h0b56dc7e;
    ram_cell[     597] = 32'hca34a464;
    ram_cell[     598] = 32'h21c54724;
    ram_cell[     599] = 32'h41e8b415;
    ram_cell[     600] = 32'he07fd9f5;
    ram_cell[     601] = 32'h2c5fb4ec;
    ram_cell[     602] = 32'h2ddb3d94;
    ram_cell[     603] = 32'h810431bf;
    ram_cell[     604] = 32'hdadd4d4a;
    ram_cell[     605] = 32'h977b2d9e;
    ram_cell[     606] = 32'h17dcd2a0;
    ram_cell[     607] = 32'hca9e596a;
    ram_cell[     608] = 32'h2e3bf718;
    ram_cell[     609] = 32'he196a4f8;
    ram_cell[     610] = 32'h8083660f;
    ram_cell[     611] = 32'h1b51de2a;
    ram_cell[     612] = 32'h72b58c71;
    ram_cell[     613] = 32'he7d78124;
    ram_cell[     614] = 32'h149d13ff;
    ram_cell[     615] = 32'h39662be0;
    ram_cell[     616] = 32'h7009debb;
    ram_cell[     617] = 32'h67d3fab5;
    ram_cell[     618] = 32'hc35a8751;
    ram_cell[     619] = 32'hcf80ae1c;
    ram_cell[     620] = 32'h69ee7b1d;
    ram_cell[     621] = 32'h076cdd22;
    ram_cell[     622] = 32'h208dd249;
    ram_cell[     623] = 32'h0f5651bf;
    ram_cell[     624] = 32'h0adc2236;
    ram_cell[     625] = 32'h9b3a0a6b;
    ram_cell[     626] = 32'hf7b7f29a;
    ram_cell[     627] = 32'h3f15b0a7;
    ram_cell[     628] = 32'hec0a1471;
    ram_cell[     629] = 32'hf426a015;
    ram_cell[     630] = 32'h3e65bc0b;
    ram_cell[     631] = 32'hc1cf7854;
    ram_cell[     632] = 32'hfec4da17;
    ram_cell[     633] = 32'h4d26e570;
    ram_cell[     634] = 32'h33d81cc4;
    ram_cell[     635] = 32'hdd3cfb76;
    ram_cell[     636] = 32'hc1bdb053;
    ram_cell[     637] = 32'h0a28fdc0;
    ram_cell[     638] = 32'h9811f39c;
    ram_cell[     639] = 32'h6ebed016;
    ram_cell[     640] = 32'h4f793bea;
    ram_cell[     641] = 32'h7e0bc11e;
    ram_cell[     642] = 32'h3a0437e7;
    ram_cell[     643] = 32'haf062b0f;
    ram_cell[     644] = 32'hd1751c64;
    ram_cell[     645] = 32'h94566e8a;
    ram_cell[     646] = 32'h3e952d28;
    ram_cell[     647] = 32'h8c00673d;
    ram_cell[     648] = 32'h309dfd0e;
    ram_cell[     649] = 32'h9264aba2;
    ram_cell[     650] = 32'h1db9c595;
    ram_cell[     651] = 32'h72d50357;
    ram_cell[     652] = 32'h2c0333c9;
    ram_cell[     653] = 32'h14b0c84d;
    ram_cell[     654] = 32'hca828cf9;
    ram_cell[     655] = 32'h8fe7355e;
    ram_cell[     656] = 32'h29bc98bd;
    ram_cell[     657] = 32'hedcde88b;
    ram_cell[     658] = 32'h090d6f7b;
    ram_cell[     659] = 32'h3f7ff0be;
    ram_cell[     660] = 32'h305a3d47;
    ram_cell[     661] = 32'h2ec5d2ed;
    ram_cell[     662] = 32'h2d609560;
    ram_cell[     663] = 32'h4c73b972;
    ram_cell[     664] = 32'hc7acef77;
    ram_cell[     665] = 32'h8216fc5e;
    ram_cell[     666] = 32'h5456b693;
    ram_cell[     667] = 32'hcbf1875d;
    ram_cell[     668] = 32'h3125b8aa;
    ram_cell[     669] = 32'hd8459251;
    ram_cell[     670] = 32'h205aa442;
    ram_cell[     671] = 32'h41526b8b;
    ram_cell[     672] = 32'h843d1f12;
    ram_cell[     673] = 32'h59f36643;
    ram_cell[     674] = 32'h0e6ec2bc;
    ram_cell[     675] = 32'h95663f4c;
    ram_cell[     676] = 32'h7f1bc6c5;
    ram_cell[     677] = 32'hff28e7d8;
    ram_cell[     678] = 32'hf8d65237;
    ram_cell[     679] = 32'h6d064c2f;
    ram_cell[     680] = 32'h04dcb7c1;
    ram_cell[     681] = 32'h630fbb97;
    ram_cell[     682] = 32'h79a1bd67;
    ram_cell[     683] = 32'h6f34c0d5;
    ram_cell[     684] = 32'h52345f0f;
    ram_cell[     685] = 32'h3fce5e6d;
    ram_cell[     686] = 32'h991d4733;
    ram_cell[     687] = 32'h9aaf437a;
    ram_cell[     688] = 32'h6983c4c7;
    ram_cell[     689] = 32'h96214e49;
    ram_cell[     690] = 32'h2d1aed2f;
    ram_cell[     691] = 32'h8774b62e;
    ram_cell[     692] = 32'h8b1580ed;
    ram_cell[     693] = 32'h39045359;
    ram_cell[     694] = 32'h376f250d;
    ram_cell[     695] = 32'he1a3b898;
    ram_cell[     696] = 32'hb5155621;
    ram_cell[     697] = 32'hc58a20cf;
    ram_cell[     698] = 32'hd03bb35c;
    ram_cell[     699] = 32'hd43e68f3;
    ram_cell[     700] = 32'h2b72994c;
    ram_cell[     701] = 32'hf717a528;
    ram_cell[     702] = 32'hf599241b;
    ram_cell[     703] = 32'hcbdb2cc4;
    ram_cell[     704] = 32'h40046e67;
    ram_cell[     705] = 32'h2aa480d7;
    ram_cell[     706] = 32'hdeec3bd4;
    ram_cell[     707] = 32'hf6916f4d;
    ram_cell[     708] = 32'h9ec5261c;
    ram_cell[     709] = 32'he597746e;
    ram_cell[     710] = 32'h4d412873;
    ram_cell[     711] = 32'h7ffb1853;
    ram_cell[     712] = 32'ha1eb1b6f;
    ram_cell[     713] = 32'h06f05b75;
    ram_cell[     714] = 32'hc38b11c1;
    ram_cell[     715] = 32'h905c7945;
    ram_cell[     716] = 32'hdb15ab8a;
    ram_cell[     717] = 32'hdf2b8f7c;
    ram_cell[     718] = 32'h038f57f0;
    ram_cell[     719] = 32'he14c82e6;
    ram_cell[     720] = 32'h8317b4f3;
    ram_cell[     721] = 32'he96b4ffa;
    ram_cell[     722] = 32'h02966a99;
    ram_cell[     723] = 32'h739a35a1;
    ram_cell[     724] = 32'hc1f7742f;
    ram_cell[     725] = 32'h8af4d0b3;
    ram_cell[     726] = 32'h42efa118;
    ram_cell[     727] = 32'hd24b92ad;
    ram_cell[     728] = 32'h4a7f9af9;
    ram_cell[     729] = 32'h901ff9db;
    ram_cell[     730] = 32'h1b10c884;
    ram_cell[     731] = 32'hbd013ca7;
    ram_cell[     732] = 32'hcdd606a4;
    ram_cell[     733] = 32'h1f423e40;
    ram_cell[     734] = 32'h6d58faa8;
    ram_cell[     735] = 32'ha66b804d;
    ram_cell[     736] = 32'hf0d72510;
    ram_cell[     737] = 32'hae97348c;
    ram_cell[     738] = 32'h52304da1;
    ram_cell[     739] = 32'h4ab83fd5;
    ram_cell[     740] = 32'h13781f4f;
    ram_cell[     741] = 32'h9385bae8;
    ram_cell[     742] = 32'h66a230f2;
    ram_cell[     743] = 32'h0644e7bb;
    ram_cell[     744] = 32'h7f7eaf64;
    ram_cell[     745] = 32'h528aaae2;
    ram_cell[     746] = 32'h7bdca174;
    ram_cell[     747] = 32'h9279af43;
    ram_cell[     748] = 32'hcd042d3e;
    ram_cell[     749] = 32'hd0ae9c1a;
    ram_cell[     750] = 32'hc8520bab;
    ram_cell[     751] = 32'h86c232f1;
    ram_cell[     752] = 32'hec4ff337;
    ram_cell[     753] = 32'h1a49574d;
    ram_cell[     754] = 32'h5070d04d;
    ram_cell[     755] = 32'h534d9ce2;
    ram_cell[     756] = 32'h29c26bc3;
    ram_cell[     757] = 32'h9bbb4e53;
    ram_cell[     758] = 32'ha53b0828;
    ram_cell[     759] = 32'h1b0fdb55;
    ram_cell[     760] = 32'h405b0154;
    ram_cell[     761] = 32'h9fa9963a;
    ram_cell[     762] = 32'h98274a6a;
    ram_cell[     763] = 32'h16fcf668;
    ram_cell[     764] = 32'hb6dfa2dd;
    ram_cell[     765] = 32'h9fb4fd8c;
    ram_cell[     766] = 32'hf8c5977b;
    ram_cell[     767] = 32'h46162c66;
end

endmodule

